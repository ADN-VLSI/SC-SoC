/////////////////////////////////////////////////////////////////////////////////////////
// Module        : Gray to Binary Code Converter
// Update at     : 19 Feb,2026
// Description   : The `gray_to_bin` module is a Gray-to-binary code converter
//                 with a data width of 8 bits.It takes an 8-bit Gray code
//                 input (`gray_i`) and converts it to its equivalent 8-bit
//                 binary output (`bin_o`).The conversion works by keeping the
//                 most significant bit (MSB) the same as the Gray code input.
//                 Each subsequent binary bit is generated by XOR-ing the
//                 previous binary bit with the current Gray code bit. This
//                 process continues from the MSB down to the least significant
//                 bit (LSB), typically implemented using a for loop to propagate
//                 the XOR operation across all 8 bits.
// Author        : Shuparna Haque (sheikhshuparna3108@gmail.com)
//
////////////////////////////////////////////////////////////////////////////////////////

module gray_2_bin #(
    // Width of the gray input and binary output
    parameter int WIDTH = 8
) (
    // Gray code input
    input  logic [WIDTH-1:0] gray_i,

    // Binary output
    output logic [WIDTH-1:0] bin_o
);

    always_comb begin
        // MSB remains the same
        bin_o[WIDTH-1] = gray_i[WIDTH-1];

        // Each lower bit is XOR of previous binary bit and current gray bit
        for (int i = WIDTH-2; i >= 0; i--) begin
            bin_o[i] = bin_o[i+1] ^ gray_i[i];
        end
    end

endmodule

                                                                               
                     
